library ieee;
use ieee.std_logic_1164.all;

--  A testbench has no ports.
entity calc_tb is
  end calc_tb;

architecture behav of calc_tb is
  --  Declaration of the component that will be instantiated.
  component calc
    port (
      op0: in std_logic;
      op1: in std_logic;
      op2: in std_logic;
      op3: in std_logic;
      op4: in std_logic;
      op5: in std_logic;
      op6: in std_logic;
      op7: in std_logic;
      clk_input: in std_logic
  ); -- output the current register content
  end component;
  --  Specifies which entity is bound with the component.
  -- for shift_reg_0: calc use entity work.calc(rtl);
  signal op0: std_logic;
  signal op1: std_logic;
  signal op2: std_logic;
  signal op3: std_logic;
  signal op4: std_logic;
  signal op5: std_logic;
  signal op6: std_logic;
  signal op7: std_logic;
  signal clk_input: std_logic;
begin
  --  Component instantiation.
  calc_0: calc
  port map (
  op0 => op0,
  op1 => op1,
  op2 => op2,
  op3 => op3,
  op4 => op4,
  op5 => op5,
  op6 => op6,
  op7 => op7,
  clk_input => clk_input
  );

  --  This process does the real job.
  process
  type pattern_type is record
    op7: std_logic;
    op6: std_logic;
    op5: std_logic;
    op4: std_logic;
    op3: std_logic;
    op2: std_logic;
    op1: std_logic;
    op0: std_logic;
    clk_input: std_logic;
  end record;
  --  The patterns to apply.
  type pattern_array is array (natural range <>) of pattern_type;
  constant patterns : pattern_array := (
  -- load $0 0
  ('1', '0', '0', '0', '0', '0', '0', '0', '1'),
  ('1', '0', '0', '0', '0', '0', '0', '0', '0'),
  -- load $1 1
  ('1', '0', '0', '1', '0', '0', '0', '1', '1'),
  ('1', '0', '0', '1', '0', '0', '0', '1', '0'),
  -- cmp1 $0 $3
  ('1', '1', '0', '0', '1', '1', '1', '1', '1'),
  ('1', '1', '0', '0', '1', '1', '1', '1', '0'),
  -- nop
  ('1', '1', '1', '1', '1', '1', '1', '1', '1'),
  ('1', '1', '1', '1', '1', '1', '1', '1', '0'),
-- nop
('1', '1', '1', '1', '1', '1', '1', '1', '1'),
('1', '1', '1', '1', '1', '1', '1', '1', '0'),
  -- prt $1 // skipped
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  -- prt $0
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),

  -- cmp1 $0 $1
  ('1', '1', '0', '0', '0', '0', '0', '1', '1'),
  ('1', '1', '0', '0', '0', '0', '0', '1', '0'),
  --nop
  ('1', '1', '1', '1', '1', '1', '1', '1', '1'),
  ('1', '1', '1', '1', '1', '1', '1', '1', '0'),
  --nop
  ('1', '1', '1', '1', '1', '1', '1', '1', '1'),
  ('1', '1', '1', '1', '1', '1', '1', '1', '0'),
  -- prt $0
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
  -- prt $1
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),

  -- load $2 2
  ('1', '0', '1', '0', '0', '0', '1', '0', '1'),
  ('1', '0', '1', '0', '0', '0', '1', '0', '0'),
  -- add $0 $1 $2
  ('0', '0', '0', '0', '0', '1', '1', '0', '1'),
  ('0', '0', '0', '0', '0', '1', '1', '0', '0'),
-- add $0 $1 $2
('0', '0', '0', '0', '0', '1', '1', '0', '1'),
('0', '0', '0', '0', '0', '1', '1', '0', '0'),
  -- load $3 3
  ('1', '0', '1', '1', '0', '0', '1', '1', '1'),
  ('1', '0', '1', '1', '0', '0', '1', '1', '0'),
-- load $3 3
('1', '0', '1', '1', '0', '0', '1', '1', '1'),
('1', '0', '1', '1', '0', '0', '1', '1', '0'),
  -- cmp1 $0 $3
  ('1', '1', '0', '0', '0', '0', '1', '1', '1'),
  ('1', '1', '0', '0', '0', '0', '1', '1', '0'),
-- cmp1 $0 $3
('1', '1', '0', '0', '0', '0', '1', '1', '1'),
('1', '1', '0', '0', '0', '0', '1', '1', '0'),
--nop
('1', '1', '1', '1', '1', '1', '1', '1', '1'),
('1', '1', '1', '1', '1', '1', '1', '1', '0'),
--nop
('1', '1', '1', '1', '1', '1', '1', '1', '1'),
('1', '1', '1', '1', '1', '1', '1', '1', '0'),
  -- prt $1
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  -- prt $0
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
  -- load $2 -2
  ('1', '0', '1', '0', '1', '1', '1', '0', '1'),
  ('1', '0', '1', '0', '1', '1', '1', '0', '0'),
  -- add $0 $1 $2
  ('0', '0', '0', '0', '0', '1', '1', '0', '1'),
  ('0', '0', '0', '0', '0', '1', '1', '0', '0'),
  ---- repeat bc hazard
('0', '0', '0', '0', '0', '1', '1', '0', '1'),
('0', '0', '0', '0', '0', '1', '1', '0', '0'),
  -- load $3 -1
  ('1', '0', '1', '1', '1', '1', '1', '1', '1'),
  ('1', '0', '1', '1', '1', '1', '1', '1', '0'),
  -- cmp1 $0 $3
  ('1', '1', '0', '0', '0', '0', '1', '1', '1'),
  ('1', '1', '0', '0', '0', '0', '1', '1', '0'),
-- repeat bc hazard
('1', '1', '0', '0', '0', '0', '1', '1', '1'),
('1', '1', '0', '0', '0', '0', '1', '1', '0'),
--nop
('1', '1', '1', '1', '1', '1', '1', '1', '1'),
('1', '1', '1', '1', '1', '1', '1', '1', '0'),
--nop
('1', '1', '1', '1', '1', '1', '1', '1', '1'),
('1', '1', '1', '1', '1', '1', '1', '1', '0'),
  -- prt $1
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  -- prt $0
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),

  -- load $1 -1
  ('1', '0', '0', '1', '1', '1', '1', '1', '1'),
  ('1', '0', '0', '1', '1', '1', '1', '1', '0'),
  -- load $3 -2
  ('1', '0', '1', '1', '1', '1', '1', '0', '1'),
  ('1', '0', '1', '1', '1', '1', '1', '0', '0'),
  -- add $0 $1 $3
  ('0', '0', '0', '0', '0', '1', '1', '1', '1'),
  ('0', '0', '0', '0', '0', '1', '1', '1', '0'),
-- add $0 $1 $3
('0', '0', '0', '0', '0', '1', '1', '1', '1'),
('0', '0', '0', '0', '0', '1', '1', '1', '0'),
  -- load $3 -3
  ('1', '0', '1', '1', '1', '1', '0', '1', '1'),
  ('1', '0', '1', '1', '1', '1', '0', '1', '0'),
  -- cmp1 $0 $3
  ('1', '1', '0', '0', '0', '0', '1', '1', '1'),
  ('1', '1', '0', '0', '0', '0', '1', '1', '0'),
-- cmp1 $0 $3
('1', '1', '0', '0', '0', '0', '1', '1', '1'),
('1', '1', '0', '0', '0', '0', '1', '1', '0'),
--nop
('1', '1', '1', '1', '1', '1', '1', '1', '1'),
('1', '1', '1', '1', '1', '1', '1', '1', '0'),
--nop
('1', '1', '1', '1', '1', '1', '1', '1', '1'),
('1', '1', '1', '1', '1', '1', '1', '1', '0'),
  -- prt $1
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  -- prt $0
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),

  --('1', '0', '0', '1', '0', '0', '0', '1', '1'),
  --('1', '0', '0', '1', '0', '0', '0', '1', '0'),
  --('1', '0', '1', '0', '0', '0', '1', '0', '1'),
  --('1', '0', '1', '0', '0', '0', '1', '0', '0'),
  --('0', '0', '0', '0', '0', '1', '1', '0', '1'),
  --('0', '0', '0', '0', '0', '1', '1', '0', '0'),
  --('1', '0', '1', '1', '0', '0', '1', '1', '1'),
  --('1', '0', '1', '1', '0', '0', '1', '1', '0'),
  --('1', '1', '0', '1', '0', '0', '1', '1', '1'),
  --('1', '1', '0', '1', '0', '0', '1', '1', '0'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '0'),
  --('1', '0', '0', '1', '0', '0', '0', '1', '1'),
  --('1', '0', '0', '1', '0', '0', '0', '1', '0'),
  --('1', '0', '1', '0', '0', '0', '1', '0', '1'),
  --('1', '0', '1', '0', '0', '0', '1', '0', '0'),
  --('0', '0', '0', '0', '0', '1', '1', '0', '1'),
  --('0', '0', '0', '0', '0', '1', '1', '0', '0'),
  --('1', '0', '1', '1', '0', '0', '1', '0', '1'),
  --('1', '0', '1', '1', '0', '0', '1', '0', '0'),
  --('1', '1', '0', '0', '0', '0', '1', '1', '1'),
  --('1', '1', '0', '0', '0', '0', '1', '1', '0'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '0'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  --('1', '0', '0', '1', '0', '0', '0', '1', '1'),
  --('1', '0', '0', '1', '0', '0', '0', '1', '0'),
  --('1', '0', '1', '0', '0', '0', '1', '0', '1'),
  --('1', '0', '1', '0', '0', '0', '1', '0', '0'),
  --('0', '0', '0', '0', '0', '1', '1', '0', '1'),
  --('0', '0', '0', '0', '0', '1', '1', '0', '0'),
  --('1', '0', '1', '1', '0', '0', '1', '0', '1'),
  --('1', '0', '1', '1', '0', '0', '1', '0', '0'),
  --('1', '1', '0', '1', '0', '0', '1', '1', '1'),
  --('1', '1', '0', '1', '0', '0', '1', '1', '0'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '0'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '0'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  --('1', '0', '0', '0', '0', '0', '0', '1', '1'),
  --('1', '0', '0', '0', '0', '0', '0', '1', '0'),
  --('1', '0', '0', '1', '0', '1', '1', '1', '1'),
  --('1', '0', '0', '1', '0', '1', '1', '1', '0'),
  --('0', '1', '0', '1', '0', '1', '0', '0', '1'),
  --('0', '1', '0', '1', '0', '1', '0', '0', '0'),
  --('1', '0', '1', '1', '0', '1', '1', '0', '1'),
  --('1', '0', '1', '1', '0', '1', '1', '0', '0'),
  --('1', '1', '0', '0', '0', '1', '1', '1', '1'),
  --('1', '1', '0', '0', '0', '1', '1', '1', '0'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '0'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  --('1', '0', '0', '0', '0', '0', '0', '1', '1'),
  --('1', '0', '0', '0', '0', '0', '0', '1', '0'),
  --('1', '0', '0', '1', '0', '1', '1', '1', '1'),
  --('1', '0', '0', '1', '0', '1', '1', '1', '0'),
  --('0', '1', '0', '1', '0', '1', '0', '0', '1'),
  --('0', '1', '0', '1', '0', '1', '0', '0', '0'),
  --('1', '0', '1', '1', '0', '1', '1', '0', '1'),
  --('1', '0', '1', '1', '0', '1', '1', '0', '0'),
  --('1', '1', '0', '1', '0', '1', '1', '1', '1'),
  --('1', '1', '0', '1', '0', '1', '1', '1', '0'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '0'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '0'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  --('1', '0', '0', '0', '0', '0', '0', '1', '1'),
  --('1', '0', '0', '0', '0', '0', '0', '1', '0'),
  --('1', '0', '0', '1', '0', '1', '1', '1', '1'),
  --('1', '0', '0', '1', '0', '1', '1', '1', '0'),
  --('0', '1', '0', '1', '0', '1', '0', '0', '1'),
  --('0', '1', '0', '1', '0', '1', '0', '0', '0'),
  --('1', '0', '1', '1', '0', '0', '1', '0', '1'),
  --('1', '0', '1', '1', '0', '0', '1', '0', '0'),
  --('1', '1', '0', '0', '0', '1', '1', '1', '1'),
  --('1', '1', '0', '0', '0', '1', '1', '1', '0'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '0'),
  --('1', '0', '0', '0', '1', '1', '1', '0', '1'),
  --('1', '0', '0', '0', '1', '1', '1', '0', '0'),
  --('1', '0', '0', '1', '1', '1', '1', '1', '1'),
  --('1', '0', '0', '1', '1', '1', '1', '1', '0'),
  --('0', '1', '0', '0', '0', '0', '0', '1', '1'),
  --('0', '1', '0', '0', '0', '0', '0', '1', '0'),
  --('1', '1', '0', '0', '0', '0', '0', '1', '1'),
  --('1', '1', '0', '0', '0', '0', '0', '1', '0'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '0'),
  --('1', '0', '0', '0', '1', '1', '1', '0', '1'),
  --('1', '0', '0', '0', '1', '1', '1', '0', '0'),
  --('1', '0', '0', '1', '0', '0', '0', '1', '1'),
  --('1', '0', '0', '1', '0', '0', '0', '1', '0'),
  --('1', '0', '1', '1', '1', '1', '0', '1', '1'),
  --('1', '0', '1', '1', '1', '1', '0', '1', '0'),
  --('0', '1', '0', '0', '0', '0', '0', '1', '1'),
  --('0', '1', '0', '0', '0', '0', '0', '1', '0'),
  --('1', '1', '0', '0', '0', '0', '1', '1', '1'),
  --('1', '1', '0', '0', '0', '0', '1', '1', '0'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '0', '0', '0', '0'),
  --('1', '0', '0', '0', '1', '0', '0', '0', '1'),
  --('1', '0', '0', '0', '1', '0', '0', '0', '0'),
  --('1', '0', '0', '1', '0', '0', '0', '1', '1'),
  --('1', '0', '0', '1', '0', '0', '0', '1', '0'),
  --('1', '0', '1', '0', '0', '0', '0', '0', '1'),
  --('1', '0', '1', '0', '0', '0', '0', '0', '0'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '1'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '0'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '1'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '0'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '1'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '0'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '1'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '0'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '1'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '0'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '1'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '0'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '1'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '0'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '1'),
  --('0', '1', '1', '0', '1', '0', '0', '1', '0'),
  --('1', '1', '0', '0', '0', '0', '1', '1', '1'),
  --('1', '1', '0', '0', '0', '0', '1', '1', '0'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '0'),
  --('1', '1', '1', '0', '1', '0', '0', '0', '1'),
  --('1', '1', '1', '0', '1', '0', '0', '0', '0'),
  ----add
  --('1', '0', '0', '1', '0', '1', '1', '1', '1'),
  --('1', '0', '0', '1', '0', '1', '1', '1', '0'),
  --('0', '0', '0', '1', '0', '1', '0', '1', '1'),
  --('0', '0', '0', '1', '0', '1', '0', '1', '0'),
  --('0', '0', '0', '1', '0', '1', '0', '1', '1'),
  --('0', '0', '0', '1', '0', '1', '0', '1', '0'),
  --('0', '0', '0', '1', '0', '1', '0', '1', '1'),
  --('0', '0', '0', '1', '0', '1', '0', '1', '0'),
  --('0', '0', '0', '1', '0', '1', '0', '1', '1'),
  --('0', '0', '0', '1', '0', '1', '0', '1', '0'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  --('1', '1', '1', '0', '0', '1', '0', '0', '0')
-- nop
('1', '1', '1', '1', '1', '1', '1', '1', '1'),
('1', '1', '1', '1', '1', '1', '1', '1', '0'),
('1', '1', '1', '1', '1', '1', '1', '1', '1'),
('1', '1', '1', '1', '1', '1', '1', '1', '0')
);
  begin
    --  Check each pattern.
    for n in patterns'range loop
      --  Set the inputs.
      op0 <= patterns(n).op0;
      op1 <= patterns(n).op1;
      op2 <= patterns(n).op2;
      op3 <= patterns(n).op3;
      op4 <= patterns(n).op4;
      op5 <= patterns(n).op5;
      op6 <= patterns(n).op6;
      op7 <= patterns(n).op7;
      clk_input <= patterns(n).clk_input;
      --  Wait for the results.
      wait for 1 ns;
      --  Check the outputs.
      --assert rd = patterns(n).rd
      --report "bad rd1 value" severity error;
      --assert clk_out = patterns(n).clk_out
      --report "bad rd2 value" severity error;
    end loop;
    assert false report "end of test" severity note;
    --  Wait forever; this will finish the simulation.
    wait;
  end process;
end behav;
