library ieee;
use ieee.std_logic_1164.all;

--  A testbench has no ports.
entity calc_tb is
  end calc_tb;

architecture behav of calc_tb is
  --  Declaration of the component that will be instantiated.
  component calc
    port (
      op0: in std_logic;
      op1: in std_logic;
      op2: in std_logic;
      op3: in std_logic;
      op4: in std_logic;
      op5: in std_logic;
      op6: in std_logic;
      op7: in std_logic;
      clk_input: in std_logic
  ); -- output the current register content
  end component;
  --  Specifies which entity is bound with the component.
  -- for shift_reg_0: calc use entity work.calc(rtl);
  signal op0: std_logic;
  signal op1: std_logic;
  signal op2: std_logic;
  signal op3: std_logic;
  signal op4: std_logic;
  signal op5: std_logic;
  signal op6: std_logic;
  signal op7: std_logic;
  signal clk_input: std_logic;
begin
  --  Component instantiation.
  calc_0: calc
  port map (
  op0 => op0,
  op1 => op1,
  op2 => op2,
  op3 => op3,
  op4 => op4,
  op5 => op5,
  op6 => op6,
  op7 => op7,
  clk_input => clk_input
  );

  --  This process does the real job.
  process
  type pattern_type is record
    op7: std_logic;
    op6: std_logic;
    op5: std_logic;
    op4: std_logic;
    op3: std_logic;
    op2: std_logic;
    op1: std_logic;
    op0: std_logic;
    clk_input: std_logic;
  end record;
  --  The patterns to apply.
  type pattern_array is array (natural range <>) of pattern_type;
  constant patterns : pattern_array := (
-- 0 one clock cycle to initialize stuff
  ('0', '0', '0', '0', '0', '0', '0', '0', '1'),
  ('0', '0', '0', '0', '0', '0', '0', '0', '0'),
-- 1 li $1 7
  ('1', '0', '0', '1', '0', '1', '1', '1', '1'),
  ('1', '0', '0', '1', '0', '1', '1', '1', '0'),
-- 2 prt $1
  ('1', '1', '1', '0', '0', '1', '0', '1', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 3 li $0 0
  ('1', '0', '0', '0', '0', '0', '0', '0', '1'),
  ('1', '0', '0', '0', '0', '0', '0', '0', '0'),
-- 4 li $1 1
  ('1', '0', '0', '1', '0', '0', '0', '1', '1'),
  ('1', '0', '0', '1', '0', '0', '0', '1', '0'),
-- 5 cmp1 $0 $3
  ('1', '1', '0', '0', '0', '0', '1', '1', '1'),
  ('1', '1', '0', '0', '0', '0', '1', '1', '0'),
-- 6 prt $1
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 7 prt $0
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 8 cmp1 $0 $1
  ('1', '1', '0', '0', '0', '0', '0', '1', '1'),
  ('1', '1', '0', '0', '0', '0', '0', '1', '0'),
-- 9
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 10
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 11
  ('1', '0', '1', '0', '0', '0', '1', '0', '1'),
  ('1', '0', '1', '0', '0', '0', '1', '0', '0'),
-- 12
  ('0', '0', '0', '0', '0', '1', '1', '0', '1'),
  ('0', '0', '0', '0', '0', '1', '1', '0', '0'),
-- 13
  ('1', '0', '1', '1', '0', '0', '1', '1', '1'),
  ('1', '0', '1', '1', '0', '0', '1', '1', '0'),
-- 14
  ('1', '1', '0', '0', '0', '0', '1', '1', '1'),
  ('1', '1', '0', '0', '0', '0', '1', '1', '0'),
-- 15
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 16
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 17
  ('1', '0', '1', '0', '1', '1', '1', '0', '1'),
  ('1', '0', '1', '0', '1', '1', '1', '0', '0'),
-- 18
  ('0', '0', '0', '0', '0', '1', '1', '0', '1'),
  ('0', '0', '0', '0', '0', '1', '1', '0', '0'),
-- 19
  ('1', '0', '1', '1', '1', '1', '1', '1', '1'),
  ('1', '0', '1', '1', '1', '1', '1', '1', '0'),
-- 20
  ('1', '1', '0', '0', '0', '0', '1', '1', '1'),
  ('1', '1', '0', '0', '0', '0', '1', '1', '0'),
-- 21
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 22
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 23
  ('1', '0', '0', '1', '1', '1', '1', '1', '1'),
  ('1', '0', '0', '1', '1', '1', '1', '1', '0'),
-- 24
  ('1', '0', '1', '1', '1', '1', '1', '0', '1'),
  ('1', '0', '1', '1', '1', '1', '1', '0', '0'),
-- 25
  ('0', '0', '0', '0', '0', '1', '1', '1', '1'),
  ('0', '0', '0', '0', '0', '1', '1', '1', '0'),
-- 26
  ('1', '0', '1', '1', '1', '1', '0', '1', '1'),
  ('1', '0', '1', '1', '1', '1', '0', '1', '0'),
-- 27
  ('1', '1', '0', '0', '0', '0', '1', '1', '1'),
  ('1', '1', '0', '0', '0', '0', '1', '1', '0'),
-- 28
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 29
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 30
  ('1', '0', '0', '1', '0', '0', '0', '1', '1'),
  ('1', '0', '0', '1', '0', '0', '0', '1', '0'),
-- 31
  ('1', '0', '1', '1', '0', '0', '1', '1', '1'),
  ('1', '0', '1', '1', '0', '0', '1', '1', '0'),
-- 32
  ('0', '0', '0', '0', '0', '1', '1', '1', '1'),
  ('0', '0', '0', '0', '0', '1', '1', '1', '0'),
-- 33
  ('1', '0', '1', '1', '0', '0', '1', '1', '1'),
  ('1', '0', '1', '1', '0', '0', '1', '1', '0'),
-- 34
  ('1', '1', '0', '1', '0', '0', '1', '1', '1'),
  ('1', '1', '0', '1', '0', '0', '1', '1', '0'),
-- 35
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 36
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 37
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 38
  ('1', '0', '0', '1', '0', '0', '0', '1', '1'),
  ('1', '0', '0', '1', '0', '0', '0', '1', '0'),
-- 39
  ('1', '0', '1', '1', '0', '0', '1', '1', '1'),
  ('1', '0', '1', '1', '0', '0', '1', '1', '0'),
-- 40
  ('0', '0', '0', '0', '0', '1', '1', '1', '1'),
  ('0', '0', '0', '0', '0', '1', '1', '1', '0'),
-- 41
  ('1', '0', '1', '1', '0', '0', '1', '1', '1'),
  ('1', '0', '1', '1', '0', '0', '1', '1', '0'),
-- 42
  ('1', '1', '0', '0', '0', '0', '1', '1', '1'),
  ('1', '1', '0', '0', '0', '0', '1', '1', '0'),
-- 43
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 44
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 45
  ('1', '0', '0', '1', '0', '0', '0', '1', '1'),
  ('1', '0', '0', '1', '0', '0', '0', '1', '0'),
-- 46
  ('1', '0', '1', '1', '0', '0', '1', '1', '1'),
  ('1', '0', '1', '1', '0', '0', '1', '1', '0'),
-- 47
  ('0', '0', '0', '0', '0', '1', '1', '1', '1'),
  ('0', '0', '0', '0', '0', '1', '1', '1', '0'),
-- 48
  ('1', '0', '1', '1', '0', '0', '1', '1', '1'),
  ('1', '0', '1', '1', '0', '0', '1', '1', '0'),
-- 49
  ('1', '1', '0', '1', '0', '0', '1', '1', '1'),
  ('1', '1', '0', '1', '0', '0', '1', '1', '0'),
-- 50
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 51
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 52
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 53
  ('1', '0', '0', '0', '0', '0', '0', '1', '1'),
  ('1', '0', '0', '0', '0', '0', '0', '1', '0'),
-- 54
  ('1', '0', '0', '1', '0', '1', '1', '1', '1'),
  ('1', '0', '0', '1', '0', '1', '1', '1', '0'),
-- 55
  ('0', '1', '0', '1', '0', '1', '0', '0', '1'),
  ('0', '1', '0', '1', '0', '1', '0', '0', '0'),
-- 56
  ('1', '0', '1', '1', '0', '1', '1', '0', '1'),
  ('1', '0', '1', '1', '0', '1', '1', '0', '0'),
-- 57
  ('1', '1', '0', '0', '0', '1', '1', '1', '1'),
  ('1', '1', '0', '0', '0', '1', '1', '1', '0'),
-- 58
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 59
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 60
  ('1', '0', '0', '0', '0', '0', '0', '1', '1'),
  ('1', '0', '0', '0', '0', '0', '0', '1', '0'),
-- 61
  ('1', '0', '0', '1', '0', '1', '1', '1', '1'),
  ('1', '0', '0', '1', '0', '1', '1', '1', '0'),
-- 62
  ('0', '1', '0', '1', '0', '1', '0', '0', '1'),
  ('0', '1', '0', '1', '0', '1', '0', '0', '0'),
-- 63
  ('1', '0', '1', '1', '0', '1', '1', '0', '1'),
  ('1', '0', '1', '1', '0', '1', '1', '0', '0'),
-- 64
  ('1', '1', '0', '1', '0', '1', '1', '1', '1'),
  ('1', '1', '0', '1', '0', '1', '1', '1', '0'),
-- 65
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 66
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 67
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 68
  ('1', '0', '0', '0', '0', '0', '0', '1', '1'),
  ('1', '0', '0', '0', '0', '0', '0', '1', '0'),
-- 69
  ('1', '0', '0', '1', '0', '1', '1', '1', '1'),
  ('1', '0', '0', '1', '0', '1', '1', '1', '0'),
-- 70
  ('0', '1', '0', '1', '0', '1', '0', '0', '1'),
  ('0', '1', '0', '1', '0', '1', '0', '0', '0'),
-- 71
  ('1', '0', '1', '1', '0', '0', '1', '0', '1'),
  ('1', '0', '1', '1', '0', '0', '1', '0', '0'),
-- 72
  ('1', '1', '0', '0', '0', '1', '1', '1', '1'),
  ('1', '1', '0', '0', '0', '1', '1', '1', '0'),
-- 73
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 74
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 75
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 76
  ('1', '0', '0', '0', '1', '1', '1', '0', '1'),
  ('1', '0', '0', '0', '1', '1', '1', '0', '0'),
-- 77
  ('1', '0', '0', '1', '1', '1', '1', '1', '1'),
  ('1', '0', '0', '1', '1', '1', '1', '1', '0'),
-- 78
  ('0', '1', '0', '0', '0', '0', '0', '1', '1'),
  ('0', '1', '0', '0', '0', '0', '0', '1', '0'),
-- 79
  ('1', '1', '0', '0', '0', '0', '0', '1', '1'),
  ('1', '1', '0', '0', '0', '0', '0', '1', '0'),
-- 80
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 81
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 82
  ('1', '0', '0', '0', '1', '1', '1', '0', '1'),
  ('1', '0', '0', '0', '1', '1', '1', '0', '0'),
-- 83
  ('1', '0', '0', '1', '0', '0', '0', '1', '1'),
  ('1', '0', '0', '1', '0', '0', '0', '1', '0'),
-- 84
  ('1', '0', '1', '1', '1', '1', '0', '1', '1'),
  ('1', '0', '1', '1', '1', '1', '0', '1', '0'),
-- 85
  ('0', '1', '0', '0', '0', '0', '0', '1', '1'),
  ('0', '1', '0', '0', '0', '0', '0', '1', '0'),
-- 86
  ('1', '1', '0', '0', '0', '0', '1', '1', '1'),
  ('1', '1', '0', '0', '0', '0', '1', '1', '0'),
-- 87
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 88
  ('1', '1', '1', '0', '0', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '0', '0', '0', '0'),
-- 89
  ('1', '0', '0', '0', '1', '0', '0', '0', '1'),
  ('1', '0', '0', '0', '1', '0', '0', '0', '0'),
-- 90
  ('1', '0', '0', '1', '0', '0', '0', '1', '1'),
  ('1', '0', '0', '1', '0', '0', '0', '1', '0'),
-- 91
  ('1', '0', '1', '1', '0', '0', '0', '0', '1'),
  ('1', '0', '1', '1', '0', '0', '0', '0', '0'),
-- 92
  ('0', '1', '1', '1', '1', '1', '0', '1', '1'),
  ('0', '1', '1', '1', '1', '1', '0', '1', '0'),
-- 93
  ('0', '1', '1', '1', '1', '1', '0', '1', '1'),
  ('0', '1', '1', '1', '1', '1', '0', '1', '0'),
-- 94
  ('0', '1', '1', '1', '1', '1', '0', '1', '1'),
  ('0', '1', '1', '1', '1', '1', '0', '1', '0'),
-- 95
  ('0', '1', '1', '1', '1', '1', '0', '1', '1'),
  ('0', '1', '1', '1', '1', '1', '0', '1', '0'),
-- 96
  ('0', '1', '1', '1', '1', '1', '0', '1', '1'),
  ('0', '1', '1', '1', '1', '1', '0', '1', '0'),
-- 97
  ('0', '1', '1', '1', '1', '1', '0', '1', '1'),
  ('0', '1', '1', '1', '1', '1', '0', '1', '0'),
-- 98
  ('0', '1', '1', '1', '1', '1', '0', '1', '1'),
  ('0', '1', '1', '1', '1', '1', '0', '1', '0'),
-- 99
  ('0', '1', '1', '1', '1', '1', '0', '1', '1'),
  ('0', '1', '1', '1', '1', '1', '0', '1', '0'),
-- 100
  ('1', '1', '0', '0', '0', '0', '1', '1', '1'),
  ('1', '1', '0', '0', '0', '0', '1', '1', '0'),
-- 101
  ('1', '1', '1', '0', '0', '1', '0', '0', '1'),
  ('1', '1', '1', '0', '0', '1', '0', '0', '0'),
-- 102 
  ('1', '1', '1', '0', '1', '0', '0', '0', '1'),
  ('1', '1', '1', '0', '1', '0', '0', '0', '0'),

('0', '0', '0', '0', '0', '0', '0', '0', '1')
);
  begin
    --  Check each pattern.
    for n in patterns'range loop
      --  Set the inputs.
      op0 <= patterns(n).op0;
      op1 <= patterns(n).op1;
      op2 <= patterns(n).op2;
      op3 <= patterns(n).op3;
      op4 <= patterns(n).op4;
      op5 <= patterns(n).op5;
      op6 <= patterns(n).op6;
      op7 <= patterns(n).op7;
      clk_input <= patterns(n).clk_input;
      --  Wait for the results.
      wait for 1 ns;
      --  Check the outputs.
      --assert rd = patterns(n).rd
      --report "bad rd1 value" severity error;
      --assert clk_out = patterns(n).clk_out
      --report "bad rd2 value" severity error;
    end loop;
    assert false report "end of test" severity note;
    --  Wait forever; this will finish the simulation.
    wait;
  end process;
end behav;
